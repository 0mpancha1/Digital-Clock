library IEEE;
use IEEE.std_logic_1164.all;
USE WORK.EE_232.ALL;

entity MODULO_6_SYNC is
port(CLK : in std_logic;
		  Q : inout std_logic_vector(3 downto 0));
end entity;



