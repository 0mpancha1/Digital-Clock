library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;


entity COUNTER_ASYNC is -- Entity declaration
	port(CLK : in std_logic; -- Clock input of the counter
		  RSTN : in std_logic; -- Active low reset input of the counter
		  Q : inout std_logic_vector(3 downto 0)); -- Output state of the counter
end entity;

architecture FUNCTIONALITY of COUNTER_ASYNC is 

begin 
	process(CLK,RSTN)
	begin
		if RSTN = '0' then
			Q <= "0000" ;
		elsif CLK'event and CLK = '1' then
			Q <= Q + '1' ;
		end if;
	end process;

end FUNCTIONALITY;

			